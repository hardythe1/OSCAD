* EESchema Netlist Version 1.1 (Spice format) creation date: Sunday 09 December 2012 03:49:27 PM IST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
U1  13 12 15 4 VPLOT8_1		
v3  9 0 5		
U6  9 11 9 7 9 6 0 1 74HC04		
R3  14 0 R		
v4  14 0 5		
U10  10 9 6 15 14 4 5 0 1 74LS109		
U7  10 9 11 13 14 12 8 0 3 15 14 12 7 9 10 1 74LS109		
R2  10 0 R		
R4  9 0 R		
R1  13 0 R		
v1  13 0 PULSE		
v2  10 0 5		

.end
