* eeschema netlist version 1.1 (spice format) creation date: sunday 09 december 2012 03:49:27 pm ist

* Plotting option vplot8_1
v3  9 0 5
* 74hc04
r3  14 0 r
v4  14 0 5
* 74ls109
* 74ls109
r2  10 0 r
r4  9 0 r
r1  13 0 r
v1  13 0 pulse(0 5 0 0 0 0.5 1)
v2  10 0 5
a1 [9] [9_in]  u6adc
a2 9_in 11_out u6
a3 [11_out] [11]  u6dac
a4 [9] [9_in]  u6adc
a5 9_in 7_out u6
a6 [7_out] [7]  u6dac
a7 [9] [9_in]  u6adc
a8 9_in 6_out u6
a9 [6_out] [6]  u6dac
.model u6 d_inverter
.model u6adc adc_bridge(in_low=0.8 in_high=2.0)
.model u6dac dac_bridge(out_low=0.25 out_high=5.0 out_undef=1.8 t_rise=0.5e-9 t_fall=0.5e-9)
a10 [9 6 15 14 10] [9_in 6_in 15_in 14_in 10_in] u10adc
a11 9_in ~6_in 15_in ~14_in ~10_in 4_out 5_out u10
a12 [4_out 5_out] [4 5]  u10dac
.model u10 d_jkff
.model u10adc adc_bridge(in_low=0.8 in_high=2.0)
.model u10dac dac_bridge(out_low=0.25 out_high=5.0 out_undef=1.8 t_rise=0.5e-9 t_fall=0.5e-9)
a13 [9 11 13 14 10] [9_in 11_in 13_in 14_in 10_in] u7adc
a14 9_in ~11_in 13_in ~14_in ~10_in 12_out 8_out u7
a15 [12_out 8_out] [12 8]  u7dac
a16 [9 7 12 14 10] [9_in 7_in 12_in 14_in 10_in] u7adc
a17 9_in ~7_in 12_in ~14_in ~10_in 15_out 3_out u7
a18 [15_out 3_out] [15 3]  u7dac
.model u7 d_jkff
.model u7adc adc_bridge(in_low=0.8 in_high=2.0)
.model u7dac dac_bridge(out_low=0.25 out_high=5.0 out_undef=1.8 t_rise=0.5e-9 t_fall=0.5e-9)

.tran  100e-03 9e-00 0e-00
.plot v(13) v(12) v(15) v(4) 
.end
