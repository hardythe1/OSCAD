* EESchema Netlist Version 1.1 (Spice format) creation date: Friday 12 April 2013 05:47:09 PM IST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
U1  3 4 1 0 VPLOT8		
V1  3 1 SINE		
R1  4 0 1000		
D3  0 3 1n4007		
D4  0 1 1n4007		
D2  1 4 1n4007		
D1  3 4 1n4007		

.end
