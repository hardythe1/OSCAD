* eeschema netlist version 1.1 (spice format) creation date: sunday 05 may 2013 04:04:48 pm ist

* Plotting option vplot8_1
v1  1 0 sine(0 5 300 0 0)
c1  3 0 1u
r1  3 1 1k

.tran  5e-03 30e-03 0e-00
.plot v(1) v(3) 
.end
